`default_nettype none
module executor(
  input  var logic clk,
  input  var logic reset,
  // handshake
  input  var logic decoder_valid,
  input  var logic executor_ready,
  output var logic executor_valid,
  input  var logic accessor_ready,
  // inputs
  input  var logic [4:0]  decoder_rd(rd),
  input  var logic [31:0] decoder_reg_rs1(decoder_reg_rs1),
  input  var logic [31:0] decoder_reg_rs2(decoder_reg_rs2),
  input  var logic [31:0] decoder_rs1(decoder_rs1),
  input  var logic [31:0] decoder_rs2(decoder_rs2),
  input  var logic [31:0] decoder_mem_addr(decoder_mem_addr),
  input  var logic        is_valid_instr(is_valid_instr),
  input  var logic        is_add(is_add),
  input  var logic        is_sub(is_sub),
  input  var logic        is_xor(is_xor),
  input  var logic        is_or(is_or),
  input  var logic        is_and(is_and),
  input  var logic        is_mul(is_mul),
  input  var logic        is_mulh(is_mulh),
  input  var logic        is_mulhu(is_mulhu),
  input  var logic        is_mulhsu(is_mulhsu),
  input  var logic        is_div(is_div),
  input  var logic        is_divu(is_divu),
  input  var logic        is_rem(is_rem),
  input  var logic        is_remu(is_remu),
  input  var logic        is_sll(is_sll),
  input  var logic        is_slt(is_slt),
  input  var logic        is_sltu(is_sltu),
  input  var logic        is_srl(is_srl),
  input  var logic        is_sra(is_sra),
  input  var logic        is_lui(is_lui),
  input  var logic        is_lb(is_lb),
  input  var logic        is_lbu(is_lbu),
  input  var logic        is_lh(is_lh),
  input  var logic        is_lhu(is_lhu),
  input  var logic        is_lw(is_lw),
  input  var logic        is_sb(is_sb),
  input  var logic        is_sh(is_sh),
  input  var logic        is_sw(is_sw),
  input  var logic        is_ecall(is_ecall),
  input  var logic        is_ebreak(is_ebreak),
  input  var logic        is_csrrw(is_csrrw),
  input  var logic        is_csrrs(is_csrrs),
  input  var logic        is_csrrc(is_csrrc),
  // forwards
  output var logic [31:0] executor_mem_addr(executor_mem_addr),
  output var logic [4:0]  executor_rd(executor_rd),
  output var logic [31:0] executor_rd_data(executor_data),
  output var logic        executor_is_lui(is_lui),
  output var logic        executor_is_lb(is_lb),
  output var logic        executor_is_lbu(is_lbu),
  output var logic        executor_is_lh(is_lh),
  output var logic        executor_is_lhu(is_lhu),
  output var logic        executor_is_lw(is_lw),
  output var logic        executor_is_sb(is_sb),
  output var logic        executor_is_sh(is_sh),
  output var logic        executor_is_sw(is_sw)
);
// handshake
// state machine
endmodule
