`default_nettype none
module accessor();

endmodule
